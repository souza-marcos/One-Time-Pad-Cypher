`ifndef __CONSTANTS_V__
`define __CONSTANTS_V__

`define KEY_SIZE 4
`define MSG_SIZE 32

`endif
