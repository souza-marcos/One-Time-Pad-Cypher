`ifndef __CONSTANTS_V__
`define __CONSTANTS_V__

`define KEY_SIZE 8     // Changing for testing
`define MSG_SIZE 64

`endif
