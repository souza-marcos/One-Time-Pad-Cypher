`ifndef __CONSTANTS_V__
`define __CONSTANTS_V__

`define KEY_SIZE 16     // Changing for testing
`define MSG_SIZE 240

`endif
