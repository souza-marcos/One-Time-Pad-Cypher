// Design:		seq
// File:		sequence_tb.v
// Description: Finite State Machine (FSM) example.
//              Sequence detectors. Mealy and Moore verions. Test bench.
// Author:		Jorge Juan-Chico <jjchico@gmail.com>
// Date: 		27-11-2010 (initial version)

/*
   Lesson 6.4: Finite State Machine (FSM) examples. Sequence detectors.

   This is a test bench for modules in 'sequence.v'. The test bench applies
   identical inputs to the Mealy and Moore versions of the sequence detector
   in order to compare the output generated by each type of machine.
 */

// In this test bench the data input is synchronous with the clock but can
// be shifted with respect to the active edge of the clock (positive edge).
// This macro controls the shift time. A value of '1' is realistic since
// synchronous inputs are expected to change right after the clock edge but
// not exactly at the same time. The XSHIFT macro can be changed to see the
// effect in the machine's behavior.
//     0: input in phase with the clock's active edge.
//  1-19: input delayed with respect to the clock's active edge
`define XSHIFT 1

`timescale 1ns / 1ps

`include "sequence.v"

// Test bench

module test ();
    reg clk = 1;    // clock
    reg reset = 0;  // reset
    reg x = 0;      // input
    wire z_mealy;   // Mealy's output
    wire z_moore;   // Moore's output

    /* 'in' vector contains a 32 bit sequence that will be applied to the
     * input. 'n' is the number of bits of the sequence and 'i' is used
     * as an index to select the bits in 'in'. */
    reg [0:31] in = 32'b00100111_00001110_10010010_01010011;
    integer n = 32;
    integer i = 0;

    // Module instantiation
    seq_mealy uut_mealy (.clk(clk), .reset(reset), .x(x), .z(z_mealy));
    seq_moore uut_moore (.clk(clk), .reset(reset), .x(x), .z(z_moore));

    // Waveform generation
    initial begin
        $dumpfile("sequence_tb.vcd");
        $dumpvars(0, test);
    end

    // Clock generator (20ns period)
    always
        #10 clk = ~clk;

    // Input sequence generator
    always @(posedge clk) begin
        // desplazamiento de la entrada respecto al reloj
        #`XSHIFT;

        x = in[i];

        // We update the index and finish if all patterns have been applied
        i = i + 1;
        if (i == n)
            $finish;
    end

    // Reset
    /* An independent process controls the 'reset' signal. We do one reset
     * at the beggining for initialization and another reset during normal
     * operation. */
    initial begin
        #5   reset = 1;
        #15  reset = 0;
        #450 reset = 1;
        #20  reset = 0;
    end
endmodule

/*
   EXERCISE

   1. Compile and simulate the design with:

        $ iverilog sequence.v sequence_tb.v
        $ vvp a.out

      and display the waveforms with gtkwave:

        $ gtkwave sequence_tb.vcd

      Visualize the input and output signals and the internal states of the
      Mealy and Moore machines.

   2. Take a look at the output waveforms and answer the following questions:

      a) Are both Mealy's and Moore's outputs identical?
      b) Is the operation of the Mealy machine correct?
      c) Is the operation of the Moore machine correct?
      d) Explain the differences observed in the outputs of both machines.

   3. Repeat the simulation for various values of the macro XSHIFT between
      0 and 19. Take a look at the changes in the output of both machines.

      a) What machine output is more affected by lack of synchronization
         between the clock and the input?
      b) What type of machine do you think will be more robust against the
         presence of inputs not synchronized with the clock?

   4. Change the input sequence ('in') and check the operation of both
      machines with the new sequence.

   5. ¿What would happen if we remove (of comment-out) the block of code
      controlling the 'reset' signal in the test bench? Try to deduce the
      result by using the machine's states table and check if your right
      with the simulation. ¿Were you right?
*/
